library verilog;
use verilog.vl_types.all;
entity top_module_vlg_check_tst is
    port(
        divisible       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end top_module_vlg_check_tst;
