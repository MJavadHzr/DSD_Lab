library verilog;
use verilog.vl_types.all;
entity top_module_vlg_sample_tst is
    port(
        A_00            : in     vl_logic;
        A_01            : in     vl_logic;
        A_02            : in     vl_logic;
        A_03            : in     vl_logic;
        A_10            : in     vl_logic;
        A_11            : in     vl_logic;
        A_12            : in     vl_logic;
        A_13            : in     vl_logic;
        A_20            : in     vl_logic;
        A_21            : in     vl_logic;
        A_22            : in     vl_logic;
        A_23            : in     vl_logic;
        A_30            : in     vl_logic;
        A_31            : in     vl_logic;
        A_32            : in     vl_logic;
        A_33            : in     vl_logic;
        div_11          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end top_module_vlg_sample_tst;
