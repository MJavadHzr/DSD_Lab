library verilog;
use verilog.vl_types.all;
entity top_module_vlg_vec_tst is
end top_module_vlg_vec_tst;
